/cad/tech/Artisan.TSMC.130/aci/sc-x/lef/tsmc13_8lm.lef